// ECE178_nios_20_1.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module ECE178_nios_20_1 (
		input  wire        clk_clk,                                            //                                         clk.clk
		output wire [7:0]  gpio_external_connection_export,                    //                    gpio_external_connection.export
		output wire [31:0] hex0_3_export,                                      //                                      hex0_3.export
		output wire [31:0] hex4_7_export,                                      //                                      hex4_7.export
		input  wire [3:0]  key_export,                                         //                                         key.export
		output wire [8:0]  ledg_export,                                        //                                        ledg.export
		output wire [17:0] ledr_export,                                        //                                        ledr.export
		input  wire        reset_reset,                                        //                                       reset.reset
		input  wire [10:0] sbus_decoder_channel_0_external_connection_export,  //  sbus_decoder_channel_0_external_connection.export
		input  wire [10:0] sbus_decoder_channel_10_external_connection_export, // sbus_decoder_channel_10_external_connection.export
		input  wire [10:0] sbus_decoder_channel_11_external_connection_export, // sbus_decoder_channel_11_external_connection.export
		input  wire [10:0] sbus_decoder_channel_12_external_connection_export, // sbus_decoder_channel_12_external_connection.export
		input  wire [10:0] sbus_decoder_channel_13_external_connection_export, // sbus_decoder_channel_13_external_connection.export
		input  wire [10:0] sbus_decoder_channel_14_external_connection_export, // sbus_decoder_channel_14_external_connection.export
		input  wire [10:0] sbus_decoder_channel_15_external_connection_export, // sbus_decoder_channel_15_external_connection.export
		input  wire [10:0] sbus_decoder_channel_1_external_connection_export,  //  sbus_decoder_channel_1_external_connection.export
		input  wire [10:0] sbus_decoder_channel_2_external_connection_export,  //  sbus_decoder_channel_2_external_connection.export
		input  wire [10:0] sbus_decoder_channel_3_external_connection_export,  //  sbus_decoder_channel_3_external_connection.export
		input  wire [10:0] sbus_decoder_channel_4_external_connection_export,  //  sbus_decoder_channel_4_external_connection.export
		input  wire [10:0] sbus_decoder_channel_5_external_connection_export,  //  sbus_decoder_channel_5_external_connection.export
		input  wire [10:0] sbus_decoder_channel_6_external_connection_export,  //  sbus_decoder_channel_6_external_connection.export
		input  wire [10:0] sbus_decoder_channel_7_external_connection_export,  //  sbus_decoder_channel_7_external_connection.export
		input  wire [10:0] sbus_decoder_channel_8_external_connection_export,  //  sbus_decoder_channel_8_external_connection.export
		input  wire [10:0] sbus_decoder_channel_9_external_connection_export,  //  sbus_decoder_channel_9_external_connection.export
		output wire [15:0] sbus_decoder_reg_0_external_connection_export,      //      sbus_decoder_reg_0_external_connection.export
		output wire [15:0] sbus_decoder_reg_10_external_connection_export,     //     sbus_decoder_reg_10_external_connection.export
		output wire [15:0] sbus_decoder_reg_1_external_connection_export,      //      sbus_decoder_reg_1_external_connection.export
		output wire [15:0] sbus_decoder_reg_2_external_connection_export,      //      sbus_decoder_reg_2_external_connection.export
		output wire [15:0] sbus_decoder_reg_3_external_connection_export,      //      sbus_decoder_reg_3_external_connection.export
		output wire [15:0] sbus_decoder_reg_4_external_connection_export,      //      sbus_decoder_reg_4_external_connection.export
		output wire [15:0] sbus_decoder_reg_5_external_connection_export,      //      sbus_decoder_reg_5_external_connection.export
		output wire [15:0] sbus_decoder_reg_6_external_connection_export,      //      sbus_decoder_reg_6_external_connection.export
		output wire [15:0] sbus_decoder_reg_7_external_connection_export,      //      sbus_decoder_reg_7_external_connection.export
		output wire [15:0] sbus_decoder_reg_8_external_connection_export,      //      sbus_decoder_reg_8_external_connection.export
		output wire [15:0] sbus_decoder_reg_9_external_connection_export,      //      sbus_decoder_reg_9_external_connection.export
		output wire [12:0] sdram_addr,                                         //                                       sdram.addr
		output wire [1:0]  sdram_ba,                                           //                                            .ba
		output wire        sdram_cas_n,                                        //                                            .cas_n
		output wire        sdram_cke,                                          //                                            .cke
		output wire        sdram_cs_n,                                         //                                            .cs_n
		inout  wire [31:0] sdram_dq,                                           //                                            .dq
		output wire [3:0]  sdram_dqm,                                          //                                            .dqm
		output wire        sdram_ras_n,                                        //                                            .ras_n
		output wire        sdram_we_n,                                         //                                            .we_n
		output wire        sdram_clk_clk,                                      //                                   sdram_clk.clk
		input  wire [17:0] switches0_17_export,                                //                                switches0_17.export
		input  wire        uart_0_external_connection_rxd,                     //                  uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd                      //                                            .txd
	);

	wire         sys_sdram_pll_0_sys_clk_clk;                                 // sys_sdram_pll_0:sys_clk_clk -> [GPIO:clk, High_Res_Timer:clk, KEYS:clk, LEDG:clk, System_Timer:clk, hex0_3:clk, hex4_7:clk, irq_mapper:clk, jtag_uart_0:clk, ledr:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, nios2_gen2_0:clk, onchip_memory2_0:clk, rst_controller:clk, rst_controller_001:clk, sbus_decoder_channel_0:clk, sbus_decoder_channel_10:clk, sbus_decoder_channel_11:clk, sbus_decoder_channel_12:clk, sbus_decoder_channel_13:clk, sbus_decoder_channel_14:clk, sbus_decoder_channel_15:clk, sbus_decoder_channel_1:clk, sbus_decoder_channel_2:clk, sbus_decoder_channel_3:clk, sbus_decoder_channel_4:clk, sbus_decoder_channel_5:clk, sbus_decoder_channel_6:clk, sbus_decoder_channel_7:clk, sbus_decoder_channel_8:clk, sbus_decoder_channel_9:clk, sbus_decoder_reg_0:clk, sbus_decoder_reg_10:clk, sbus_decoder_reg_1:clk, sbus_decoder_reg_2:clk, sbus_decoder_reg_3:clk, sbus_decoder_reg_4:clk, sbus_decoder_reg_5:clk, sbus_decoder_reg_6:clk, sbus_decoder_reg_7:clk, sbus_decoder_reg_8:clk, sbus_decoder_reg_9:clk, sdram_0:clk, switches0_17:clk, uart_0:clk]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> [LEDG:reset_n, mm_interconnect_0:LEDG_reset_reset_bridge_in_reset_reset, rst_controller_001:reset_in0]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_hex0_3_s1_chipselect;                      // mm_interconnect_0:hex0_3_s1_chipselect -> hex0_3:chipselect
	wire  [31:0] mm_interconnect_0_hex0_3_s1_readdata;                        // hex0_3:readdata -> mm_interconnect_0:hex0_3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex0_3_s1_address;                         // mm_interconnect_0:hex0_3_s1_address -> hex0_3:address
	wire         mm_interconnect_0_hex0_3_s1_write;                           // mm_interconnect_0:hex0_3_s1_write -> hex0_3:write_n
	wire  [31:0] mm_interconnect_0_hex0_3_s1_writedata;                       // mm_interconnect_0:hex0_3_s1_writedata -> hex0_3:writedata
	wire         mm_interconnect_0_hex4_7_s1_chipselect;                      // mm_interconnect_0:hex4_7_s1_chipselect -> hex4_7:chipselect
	wire  [31:0] mm_interconnect_0_hex4_7_s1_readdata;                        // hex4_7:readdata -> mm_interconnect_0:hex4_7_s1_readdata
	wire   [1:0] mm_interconnect_0_hex4_7_s1_address;                         // mm_interconnect_0:hex4_7_s1_address -> hex4_7:address
	wire         mm_interconnect_0_hex4_7_s1_write;                           // mm_interconnect_0:hex4_7_s1_write -> hex4_7:write_n
	wire  [31:0] mm_interconnect_0_hex4_7_s1_writedata;                       // mm_interconnect_0:hex4_7_s1_writedata -> hex4_7:writedata
	wire  [31:0] mm_interconnect_0_switches0_17_s1_readdata;                  // switches0_17:readdata -> mm_interconnect_0:switches0_17_s1_readdata
	wire   [1:0] mm_interconnect_0_switches0_17_s1_address;                   // mm_interconnect_0:switches0_17_s1_address -> switches0_17:address
	wire         mm_interconnect_0_ledr_s1_chipselect;                        // mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                          // ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                           // mm_interconnect_0:ledr_s1_address -> ledr:address
	wire         mm_interconnect_0_ledr_s1_write;                             // mm_interconnect_0:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                         // mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	wire         mm_interconnect_0_high_res_timer_s1_chipselect;              // mm_interconnect_0:High_Res_Timer_s1_chipselect -> High_Res_Timer:chipselect
	wire  [15:0] mm_interconnect_0_high_res_timer_s1_readdata;                // High_Res_Timer:readdata -> mm_interconnect_0:High_Res_Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_high_res_timer_s1_address;                 // mm_interconnect_0:High_Res_Timer_s1_address -> High_Res_Timer:address
	wire         mm_interconnect_0_high_res_timer_s1_write;                   // mm_interconnect_0:High_Res_Timer_s1_write -> High_Res_Timer:write_n
	wire  [15:0] mm_interconnect_0_high_res_timer_s1_writedata;               // mm_interconnect_0:High_Res_Timer_s1_writedata -> High_Res_Timer:writedata
	wire         mm_interconnect_0_system_timer_s1_chipselect;                // mm_interconnect_0:System_Timer_s1_chipselect -> System_Timer:chipselect
	wire  [15:0] mm_interconnect_0_system_timer_s1_readdata;                  // System_Timer:readdata -> mm_interconnect_0:System_Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_system_timer_s1_address;                   // mm_interconnect_0:System_Timer_s1_address -> System_Timer:address
	wire         mm_interconnect_0_system_timer_s1_write;                     // mm_interconnect_0:System_Timer_s1_write -> System_Timer:write_n
	wire  [15:0] mm_interconnect_0_system_timer_s1_writedata;                 // mm_interconnect_0:System_Timer_s1_writedata -> System_Timer:writedata
	wire         mm_interconnect_0_sdram_0_s1_chipselect;                     // mm_interconnect_0:sdram_0_s1_chipselect -> sdram_0:az_cs
	wire  [31:0] mm_interconnect_0_sdram_0_s1_readdata;                       // sdram_0:za_data -> mm_interconnect_0:sdram_0_s1_readdata
	wire         mm_interconnect_0_sdram_0_s1_waitrequest;                    // sdram_0:za_waitrequest -> mm_interconnect_0:sdram_0_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_0_s1_address;                        // mm_interconnect_0:sdram_0_s1_address -> sdram_0:az_addr
	wire         mm_interconnect_0_sdram_0_s1_read;                           // mm_interconnect_0:sdram_0_s1_read -> sdram_0:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_0_s1_byteenable;                     // mm_interconnect_0:sdram_0_s1_byteenable -> sdram_0:az_be_n
	wire         mm_interconnect_0_sdram_0_s1_readdatavalid;                  // sdram_0:za_valid -> mm_interconnect_0:sdram_0_s1_readdatavalid
	wire         mm_interconnect_0_sdram_0_s1_write;                          // mm_interconnect_0:sdram_0_s1_write -> sdram_0:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_0_s1_writedata;                      // mm_interconnect_0:sdram_0_s1_writedata -> sdram_0:az_data
	wire         mm_interconnect_0_ledg_s1_chipselect;                        // mm_interconnect_0:LEDG_s1_chipselect -> LEDG:chipselect
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                          // LEDG:readdata -> mm_interconnect_0:LEDG_s1_readdata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                           // mm_interconnect_0:LEDG_s1_address -> LEDG:address
	wire         mm_interconnect_0_ledg_s1_write;                             // mm_interconnect_0:LEDG_s1_write -> LEDG:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                         // mm_interconnect_0:LEDG_s1_writedata -> LEDG:writedata
	wire         mm_interconnect_0_keys_s1_chipselect;                        // mm_interconnect_0:KEYS_s1_chipselect -> KEYS:chipselect
	wire  [31:0] mm_interconnect_0_keys_s1_readdata;                          // KEYS:readdata -> mm_interconnect_0:KEYS_s1_readdata
	wire   [1:0] mm_interconnect_0_keys_s1_address;                           // mm_interconnect_0:KEYS_s1_address -> KEYS:address
	wire         mm_interconnect_0_keys_s1_write;                             // mm_interconnect_0:KEYS_s1_write -> KEYS:write_n
	wire  [31:0] mm_interconnect_0_keys_s1_writedata;                         // mm_interconnect_0:KEYS_s1_writedata -> KEYS:writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;                      // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                        // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                         // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                            // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                   // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                           // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                       // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         mm_interconnect_0_gpio_s1_chipselect;                        // mm_interconnect_0:GPIO_s1_chipselect -> GPIO:chipselect
	wire  [31:0] mm_interconnect_0_gpio_s1_readdata;                          // GPIO:readdata -> mm_interconnect_0:GPIO_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio_s1_address;                           // mm_interconnect_0:GPIO_s1_address -> GPIO:address
	wire         mm_interconnect_0_gpio_s1_write;                             // mm_interconnect_0:GPIO_s1_write -> GPIO:write_n
	wire  [31:0] mm_interconnect_0_gpio_s1_writedata;                         // mm_interconnect_0:GPIO_s1_writedata -> GPIO:writedata
	wire         mm_interconnect_0_sbus_decoder_reg_0_s1_chipselect;          // mm_interconnect_0:sbus_decoder_reg_0_s1_chipselect -> sbus_decoder_reg_0:chipselect
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_0_s1_readdata;            // sbus_decoder_reg_0:readdata -> mm_interconnect_0:sbus_decoder_reg_0_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_reg_0_s1_address;             // mm_interconnect_0:sbus_decoder_reg_0_s1_address -> sbus_decoder_reg_0:address
	wire         mm_interconnect_0_sbus_decoder_reg_0_s1_write;               // mm_interconnect_0:sbus_decoder_reg_0_s1_write -> sbus_decoder_reg_0:write_n
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_0_s1_writedata;           // mm_interconnect_0:sbus_decoder_reg_0_s1_writedata -> sbus_decoder_reg_0:writedata
	wire         mm_interconnect_0_sbus_decoder_reg_1_s1_chipselect;          // mm_interconnect_0:sbus_decoder_reg_1_s1_chipselect -> sbus_decoder_reg_1:chipselect
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_1_s1_readdata;            // sbus_decoder_reg_1:readdata -> mm_interconnect_0:sbus_decoder_reg_1_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_reg_1_s1_address;             // mm_interconnect_0:sbus_decoder_reg_1_s1_address -> sbus_decoder_reg_1:address
	wire         mm_interconnect_0_sbus_decoder_reg_1_s1_write;               // mm_interconnect_0:sbus_decoder_reg_1_s1_write -> sbus_decoder_reg_1:write_n
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_1_s1_writedata;           // mm_interconnect_0:sbus_decoder_reg_1_s1_writedata -> sbus_decoder_reg_1:writedata
	wire         mm_interconnect_0_sbus_decoder_reg_2_s1_chipselect;          // mm_interconnect_0:sbus_decoder_reg_2_s1_chipselect -> sbus_decoder_reg_2:chipselect
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_2_s1_readdata;            // sbus_decoder_reg_2:readdata -> mm_interconnect_0:sbus_decoder_reg_2_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_reg_2_s1_address;             // mm_interconnect_0:sbus_decoder_reg_2_s1_address -> sbus_decoder_reg_2:address
	wire         mm_interconnect_0_sbus_decoder_reg_2_s1_write;               // mm_interconnect_0:sbus_decoder_reg_2_s1_write -> sbus_decoder_reg_2:write_n
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_2_s1_writedata;           // mm_interconnect_0:sbus_decoder_reg_2_s1_writedata -> sbus_decoder_reg_2:writedata
	wire         mm_interconnect_0_sbus_decoder_reg_3_s1_chipselect;          // mm_interconnect_0:sbus_decoder_reg_3_s1_chipselect -> sbus_decoder_reg_3:chipselect
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_3_s1_readdata;            // sbus_decoder_reg_3:readdata -> mm_interconnect_0:sbus_decoder_reg_3_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_reg_3_s1_address;             // mm_interconnect_0:sbus_decoder_reg_3_s1_address -> sbus_decoder_reg_3:address
	wire         mm_interconnect_0_sbus_decoder_reg_3_s1_write;               // mm_interconnect_0:sbus_decoder_reg_3_s1_write -> sbus_decoder_reg_3:write_n
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_3_s1_writedata;           // mm_interconnect_0:sbus_decoder_reg_3_s1_writedata -> sbus_decoder_reg_3:writedata
	wire         mm_interconnect_0_sbus_decoder_reg_4_s1_chipselect;          // mm_interconnect_0:sbus_decoder_reg_4_s1_chipselect -> sbus_decoder_reg_4:chipselect
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_4_s1_readdata;            // sbus_decoder_reg_4:readdata -> mm_interconnect_0:sbus_decoder_reg_4_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_reg_4_s1_address;             // mm_interconnect_0:sbus_decoder_reg_4_s1_address -> sbus_decoder_reg_4:address
	wire         mm_interconnect_0_sbus_decoder_reg_4_s1_write;               // mm_interconnect_0:sbus_decoder_reg_4_s1_write -> sbus_decoder_reg_4:write_n
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_4_s1_writedata;           // mm_interconnect_0:sbus_decoder_reg_4_s1_writedata -> sbus_decoder_reg_4:writedata
	wire         mm_interconnect_0_sbus_decoder_reg_5_s1_chipselect;          // mm_interconnect_0:sbus_decoder_reg_5_s1_chipselect -> sbus_decoder_reg_5:chipselect
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_5_s1_readdata;            // sbus_decoder_reg_5:readdata -> mm_interconnect_0:sbus_decoder_reg_5_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_reg_5_s1_address;             // mm_interconnect_0:sbus_decoder_reg_5_s1_address -> sbus_decoder_reg_5:address
	wire         mm_interconnect_0_sbus_decoder_reg_5_s1_write;               // mm_interconnect_0:sbus_decoder_reg_5_s1_write -> sbus_decoder_reg_5:write_n
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_5_s1_writedata;           // mm_interconnect_0:sbus_decoder_reg_5_s1_writedata -> sbus_decoder_reg_5:writedata
	wire         mm_interconnect_0_sbus_decoder_reg_6_s1_chipselect;          // mm_interconnect_0:sbus_decoder_reg_6_s1_chipselect -> sbus_decoder_reg_6:chipselect
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_6_s1_readdata;            // sbus_decoder_reg_6:readdata -> mm_interconnect_0:sbus_decoder_reg_6_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_reg_6_s1_address;             // mm_interconnect_0:sbus_decoder_reg_6_s1_address -> sbus_decoder_reg_6:address
	wire         mm_interconnect_0_sbus_decoder_reg_6_s1_write;               // mm_interconnect_0:sbus_decoder_reg_6_s1_write -> sbus_decoder_reg_6:write_n
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_6_s1_writedata;           // mm_interconnect_0:sbus_decoder_reg_6_s1_writedata -> sbus_decoder_reg_6:writedata
	wire         mm_interconnect_0_sbus_decoder_reg_7_s1_chipselect;          // mm_interconnect_0:sbus_decoder_reg_7_s1_chipselect -> sbus_decoder_reg_7:chipselect
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_7_s1_readdata;            // sbus_decoder_reg_7:readdata -> mm_interconnect_0:sbus_decoder_reg_7_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_reg_7_s1_address;             // mm_interconnect_0:sbus_decoder_reg_7_s1_address -> sbus_decoder_reg_7:address
	wire         mm_interconnect_0_sbus_decoder_reg_7_s1_write;               // mm_interconnect_0:sbus_decoder_reg_7_s1_write -> sbus_decoder_reg_7:write_n
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_7_s1_writedata;           // mm_interconnect_0:sbus_decoder_reg_7_s1_writedata -> sbus_decoder_reg_7:writedata
	wire         mm_interconnect_0_sbus_decoder_reg_8_s1_chipselect;          // mm_interconnect_0:sbus_decoder_reg_8_s1_chipselect -> sbus_decoder_reg_8:chipselect
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_8_s1_readdata;            // sbus_decoder_reg_8:readdata -> mm_interconnect_0:sbus_decoder_reg_8_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_reg_8_s1_address;             // mm_interconnect_0:sbus_decoder_reg_8_s1_address -> sbus_decoder_reg_8:address
	wire         mm_interconnect_0_sbus_decoder_reg_8_s1_write;               // mm_interconnect_0:sbus_decoder_reg_8_s1_write -> sbus_decoder_reg_8:write_n
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_8_s1_writedata;           // mm_interconnect_0:sbus_decoder_reg_8_s1_writedata -> sbus_decoder_reg_8:writedata
	wire         mm_interconnect_0_sbus_decoder_reg_9_s1_chipselect;          // mm_interconnect_0:sbus_decoder_reg_9_s1_chipselect -> sbus_decoder_reg_9:chipselect
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_9_s1_readdata;            // sbus_decoder_reg_9:readdata -> mm_interconnect_0:sbus_decoder_reg_9_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_reg_9_s1_address;             // mm_interconnect_0:sbus_decoder_reg_9_s1_address -> sbus_decoder_reg_9:address
	wire         mm_interconnect_0_sbus_decoder_reg_9_s1_write;               // mm_interconnect_0:sbus_decoder_reg_9_s1_write -> sbus_decoder_reg_9:write_n
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_9_s1_writedata;           // mm_interconnect_0:sbus_decoder_reg_9_s1_writedata -> sbus_decoder_reg_9:writedata
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_0_s1_readdata;        // sbus_decoder_channel_0:readdata -> mm_interconnect_0:sbus_decoder_channel_0_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_0_s1_address;         // mm_interconnect_0:sbus_decoder_channel_0_s1_address -> sbus_decoder_channel_0:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_1_s1_readdata;        // sbus_decoder_channel_1:readdata -> mm_interconnect_0:sbus_decoder_channel_1_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_1_s1_address;         // mm_interconnect_0:sbus_decoder_channel_1_s1_address -> sbus_decoder_channel_1:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_2_s1_readdata;        // sbus_decoder_channel_2:readdata -> mm_interconnect_0:sbus_decoder_channel_2_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_2_s1_address;         // mm_interconnect_0:sbus_decoder_channel_2_s1_address -> sbus_decoder_channel_2:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_3_s1_readdata;        // sbus_decoder_channel_3:readdata -> mm_interconnect_0:sbus_decoder_channel_3_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_3_s1_address;         // mm_interconnect_0:sbus_decoder_channel_3_s1_address -> sbus_decoder_channel_3:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_4_s1_readdata;        // sbus_decoder_channel_4:readdata -> mm_interconnect_0:sbus_decoder_channel_4_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_4_s1_address;         // mm_interconnect_0:sbus_decoder_channel_4_s1_address -> sbus_decoder_channel_4:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_5_s1_readdata;        // sbus_decoder_channel_5:readdata -> mm_interconnect_0:sbus_decoder_channel_5_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_5_s1_address;         // mm_interconnect_0:sbus_decoder_channel_5_s1_address -> sbus_decoder_channel_5:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_6_s1_readdata;        // sbus_decoder_channel_6:readdata -> mm_interconnect_0:sbus_decoder_channel_6_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_6_s1_address;         // mm_interconnect_0:sbus_decoder_channel_6_s1_address -> sbus_decoder_channel_6:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_7_s1_readdata;        // sbus_decoder_channel_7:readdata -> mm_interconnect_0:sbus_decoder_channel_7_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_7_s1_address;         // mm_interconnect_0:sbus_decoder_channel_7_s1_address -> sbus_decoder_channel_7:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_8_s1_readdata;        // sbus_decoder_channel_8:readdata -> mm_interconnect_0:sbus_decoder_channel_8_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_8_s1_address;         // mm_interconnect_0:sbus_decoder_channel_8_s1_address -> sbus_decoder_channel_8:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_9_s1_readdata;        // sbus_decoder_channel_9:readdata -> mm_interconnect_0:sbus_decoder_channel_9_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_9_s1_address;         // mm_interconnect_0:sbus_decoder_channel_9_s1_address -> sbus_decoder_channel_9:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_10_s1_readdata;       // sbus_decoder_channel_10:readdata -> mm_interconnect_0:sbus_decoder_channel_10_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_10_s1_address;        // mm_interconnect_0:sbus_decoder_channel_10_s1_address -> sbus_decoder_channel_10:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_11_s1_readdata;       // sbus_decoder_channel_11:readdata -> mm_interconnect_0:sbus_decoder_channel_11_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_11_s1_address;        // mm_interconnect_0:sbus_decoder_channel_11_s1_address -> sbus_decoder_channel_11:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_12_s1_readdata;       // sbus_decoder_channel_12:readdata -> mm_interconnect_0:sbus_decoder_channel_12_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_12_s1_address;        // mm_interconnect_0:sbus_decoder_channel_12_s1_address -> sbus_decoder_channel_12:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_13_s1_readdata;       // sbus_decoder_channel_13:readdata -> mm_interconnect_0:sbus_decoder_channel_13_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_13_s1_address;        // mm_interconnect_0:sbus_decoder_channel_13_s1_address -> sbus_decoder_channel_13:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_14_s1_readdata;       // sbus_decoder_channel_14:readdata -> mm_interconnect_0:sbus_decoder_channel_14_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_14_s1_address;        // mm_interconnect_0:sbus_decoder_channel_14_s1_address -> sbus_decoder_channel_14:address
	wire  [31:0] mm_interconnect_0_sbus_decoder_channel_15_s1_readdata;       // sbus_decoder_channel_15:readdata -> mm_interconnect_0:sbus_decoder_channel_15_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_channel_15_s1_address;        // mm_interconnect_0:sbus_decoder_channel_15_s1_address -> sbus_decoder_channel_15:address
	wire         mm_interconnect_0_sbus_decoder_reg_10_s1_chipselect;         // mm_interconnect_0:sbus_decoder_reg_10_s1_chipselect -> sbus_decoder_reg_10:chipselect
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_10_s1_readdata;           // sbus_decoder_reg_10:readdata -> mm_interconnect_0:sbus_decoder_reg_10_s1_readdata
	wire   [1:0] mm_interconnect_0_sbus_decoder_reg_10_s1_address;            // mm_interconnect_0:sbus_decoder_reg_10_s1_address -> sbus_decoder_reg_10:address
	wire         mm_interconnect_0_sbus_decoder_reg_10_s1_write;              // mm_interconnect_0:sbus_decoder_reg_10_s1_write -> sbus_decoder_reg_10:write_n
	wire  [31:0] mm_interconnect_0_sbus_decoder_reg_10_s1_writedata;          // mm_interconnect_0:sbus_decoder_reg_10_s1_writedata -> sbus_decoder_reg_10:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // High_Res_Timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // System_Timer:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // KEYS:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                    // uart_0:irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [GPIO:reset_n, mm_interconnect_0:uart_0_reset_reset_bridge_in_reset_reset, sbus_decoder_channel_0:reset_n, sbus_decoder_channel_10:reset_n, sbus_decoder_channel_11:reset_n, sbus_decoder_channel_12:reset_n, sbus_decoder_channel_13:reset_n, sbus_decoder_channel_14:reset_n, sbus_decoder_channel_15:reset_n, sbus_decoder_channel_1:reset_n, sbus_decoder_channel_2:reset_n, sbus_decoder_channel_3:reset_n, sbus_decoder_channel_4:reset_n, sbus_decoder_channel_5:reset_n, sbus_decoder_channel_6:reset_n, sbus_decoder_channel_7:reset_n, sbus_decoder_channel_8:reset_n, sbus_decoder_channel_9:reset_n, sbus_decoder_reg_0:reset_n, sbus_decoder_reg_10:reset_n, sbus_decoder_reg_1:reset_n, sbus_decoder_reg_2:reset_n, sbus_decoder_reg_3:reset_n, sbus_decoder_reg_4:reset_n, sbus_decoder_reg_5:reset_n, sbus_decoder_reg_6:reset_n, sbus_decoder_reg_7:reset_n, sbus_decoder_reg_8:reset_n, sbus_decoder_reg_9:reset_n, uart_0:reset_n]
	wire         sys_sdram_pll_0_reset_source_reset;                          // sys_sdram_pll_0:reset_source_reset -> [rst_controller:reset_in0, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [High_Res_Timer:reset_n, KEYS:reset_n, System_Timer:reset_n, hex0_3:reset_n, hex4_7:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, ledr:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sdram_0:reset_n, switches0_17:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	ECE178_nios_20_1_GPIO gpio (
		.clk        (sys_sdram_pll_0_sys_clk_clk),          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio_s1_readdata),   //                    .readdata
		.out_port   (gpio_external_connection_export)       // external_connection.export
	);

	ECE178_nios_20_1_High_Res_Timer high_res_timer (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                    //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),            // reset.reset_n
		.address    (mm_interconnect_0_high_res_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_high_res_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_high_res_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_high_res_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_high_res_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                        //   irq.irq
	);

	ECE178_nios_20_1_KEYS keys (
		.clk        (sys_sdram_pll_0_sys_clk_clk),          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_keys_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keys_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keys_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keys_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keys_s1_readdata),   //                    .readdata
		.in_port    (key_export),                           // external_connection.export
		.irq        (irq_mapper_receiver3_irq)              //                 irq.irq
	);

	ECE178_nios_20_1_LEDG ledg (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //                 clk.clk
		.reset_n    (~nios2_gen2_0_debug_reset_request_reset), //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),       //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),        //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),     //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect),    //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),      //                    .readdata
		.out_port   (ledg_export)                              // external_connection.export
	);

	ECE178_nios_20_1_System_Timer system_timer (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                  //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_system_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_system_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_system_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_system_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_system_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                      //   irq.irq
	);

	ECE178_nios_20_1_hex0_3 hex0_3 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_hex0_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex0_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex0_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex0_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex0_3_s1_readdata),   //                    .readdata
		.out_port   (hex0_3_export)                           // external_connection.export
	);

	ECE178_nios_20_1_hex0_3 hex4_7 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_hex4_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex4_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex4_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex4_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex4_7_s1_readdata),   //                    .readdata
		.out_port   (hex4_7_export)                           // external_connection.export
	);

	ECE178_nios_20_1_jtag_uart_0 jtag_uart_0 (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                                 //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	ECE178_nios_20_1_ledr ledr (
		.clk        (sys_sdram_pll_0_sys_clk_clk),          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	ECE178_nios_20_1_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (sys_sdram_pll_0_sys_clk_clk),                                //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	ECE178_nios_20_1_onchip_memory2_0 onchip_memory2_0 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                      //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_0 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_0_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_0_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_1 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_1_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_1_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_10 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_10_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_10_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_10_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_11 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_11_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_11_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_11_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_12 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_12_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_12_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_12_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_13 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_13_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_13_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_13_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_14 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_14_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_14_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_14_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_15 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_15_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_15_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_15_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_2 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_2_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_2_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_3 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_3_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_3_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_4 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_4_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_4_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_5 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_5_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_5_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_5_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_6 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_6_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_6_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_6_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_7 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_7_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_7_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_7_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_8 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_8_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_8_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_8_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_channel_0 sbus_decoder_channel_9 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address  (mm_interconnect_0_sbus_decoder_channel_9_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sbus_decoder_channel_9_s1_readdata), //                    .readdata
		.in_port  (sbus_decoder_channel_9_external_connection_export)     // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_reg_0 sbus_decoder_reg_0 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_sbus_decoder_reg_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sbus_decoder_reg_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sbus_decoder_reg_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sbus_decoder_reg_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sbus_decoder_reg_0_s1_readdata),   //                    .readdata
		.out_port   (sbus_decoder_reg_0_external_connection_export)       // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_reg_0 sbus_decoder_reg_1 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_sbus_decoder_reg_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sbus_decoder_reg_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sbus_decoder_reg_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sbus_decoder_reg_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sbus_decoder_reg_1_s1_readdata),   //                    .readdata
		.out_port   (sbus_decoder_reg_1_external_connection_export)       // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_reg_0 sbus_decoder_reg_10 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (mm_interconnect_0_sbus_decoder_reg_10_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sbus_decoder_reg_10_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sbus_decoder_reg_10_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sbus_decoder_reg_10_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sbus_decoder_reg_10_s1_readdata),   //                    .readdata
		.out_port   (sbus_decoder_reg_10_external_connection_export)       // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_reg_0 sbus_decoder_reg_2 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_sbus_decoder_reg_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sbus_decoder_reg_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sbus_decoder_reg_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sbus_decoder_reg_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sbus_decoder_reg_2_s1_readdata),   //                    .readdata
		.out_port   (sbus_decoder_reg_2_external_connection_export)       // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_reg_0 sbus_decoder_reg_3 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_sbus_decoder_reg_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sbus_decoder_reg_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sbus_decoder_reg_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sbus_decoder_reg_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sbus_decoder_reg_3_s1_readdata),   //                    .readdata
		.out_port   (sbus_decoder_reg_3_external_connection_export)       // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_reg_0 sbus_decoder_reg_4 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_sbus_decoder_reg_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sbus_decoder_reg_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sbus_decoder_reg_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sbus_decoder_reg_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sbus_decoder_reg_4_s1_readdata),   //                    .readdata
		.out_port   (sbus_decoder_reg_4_external_connection_export)       // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_reg_0 sbus_decoder_reg_5 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_sbus_decoder_reg_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sbus_decoder_reg_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sbus_decoder_reg_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sbus_decoder_reg_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sbus_decoder_reg_5_s1_readdata),   //                    .readdata
		.out_port   (sbus_decoder_reg_5_external_connection_export)       // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_reg_0 sbus_decoder_reg_6 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_sbus_decoder_reg_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sbus_decoder_reg_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sbus_decoder_reg_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sbus_decoder_reg_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sbus_decoder_reg_6_s1_readdata),   //                    .readdata
		.out_port   (sbus_decoder_reg_6_external_connection_export)       // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_reg_0 sbus_decoder_reg_7 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_sbus_decoder_reg_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sbus_decoder_reg_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sbus_decoder_reg_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sbus_decoder_reg_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sbus_decoder_reg_7_s1_readdata),   //                    .readdata
		.out_port   (sbus_decoder_reg_7_external_connection_export)       // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_reg_0 sbus_decoder_reg_8 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_sbus_decoder_reg_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sbus_decoder_reg_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sbus_decoder_reg_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sbus_decoder_reg_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sbus_decoder_reg_8_s1_readdata),   //                    .readdata
		.out_port   (sbus_decoder_reg_8_external_connection_export)       // external_connection.export
	);

	ECE178_nios_20_1_sbus_decoder_reg_0 sbus_decoder_reg_9 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_sbus_decoder_reg_9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sbus_decoder_reg_9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sbus_decoder_reg_9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sbus_decoder_reg_9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sbus_decoder_reg_9_s1_readdata),   //                    .readdata
		.out_port   (sbus_decoder_reg_9_external_connection_export)       // external_connection.export
	);

	ECE178_nios_20_1_sdram_0 sdram_0 (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),        // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                 //  wire.export
		.zs_ba          (sdram_ba),                                   //      .export
		.zs_cas_n       (sdram_cas_n),                                //      .export
		.zs_cke         (sdram_cke),                                  //      .export
		.zs_cs_n        (sdram_cs_n),                                 //      .export
		.zs_dq          (sdram_dq),                                   //      .export
		.zs_dqm         (sdram_dqm),                                  //      .export
		.zs_ras_n       (sdram_ras_n),                                //      .export
		.zs_we_n        (sdram_we_n)                                  //      .export
	);

	ECE178_nios_20_1_switches0_17 switches0_17 (
		.clk      (sys_sdram_pll_0_sys_clk_clk),                //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches0_17_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches0_17_s1_readdata), //                    .readdata
		.in_port  (switches0_17_export)                         // external_connection.export
	);

	ECE178_nios_20_1_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (reset_reset),                        //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_0_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset (sys_sdram_pll_0_reset_source_reset)  // reset_source.reset
	);

	ECE178_nios_20_1_uart_0 uart_0 (
		.clk           (sys_sdram_pll_0_sys_clk_clk),               //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_0_external_connection_rxd),            // external_connection.export
		.txd           (uart_0_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver4_irq)                   //                 irq.irq
	);

	ECE178_nios_20_1_mm_interconnect_0 mm_interconnect_0 (
		.sys_sdram_pll_0_sys_clk_clk                    (sys_sdram_pll_0_sys_clk_clk),                                 //                  sys_sdram_pll_0_sys_clk.clk
		.LEDG_reset_reset_bridge_in_reset_reset         (nios2_gen2_0_debug_reset_request_reset),                      //         LEDG_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.uart_0_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                              //       uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.GPIO_s1_address                                (mm_interconnect_0_gpio_s1_address),                           //                                  GPIO_s1.address
		.GPIO_s1_write                                  (mm_interconnect_0_gpio_s1_write),                             //                                         .write
		.GPIO_s1_readdata                               (mm_interconnect_0_gpio_s1_readdata),                          //                                         .readdata
		.GPIO_s1_writedata                              (mm_interconnect_0_gpio_s1_writedata),                         //                                         .writedata
		.GPIO_s1_chipselect                             (mm_interconnect_0_gpio_s1_chipselect),                        //                                         .chipselect
		.hex0_3_s1_address                              (mm_interconnect_0_hex0_3_s1_address),                         //                                hex0_3_s1.address
		.hex0_3_s1_write                                (mm_interconnect_0_hex0_3_s1_write),                           //                                         .write
		.hex0_3_s1_readdata                             (mm_interconnect_0_hex0_3_s1_readdata),                        //                                         .readdata
		.hex0_3_s1_writedata                            (mm_interconnect_0_hex0_3_s1_writedata),                       //                                         .writedata
		.hex0_3_s1_chipselect                           (mm_interconnect_0_hex0_3_s1_chipselect),                      //                                         .chipselect
		.hex4_7_s1_address                              (mm_interconnect_0_hex4_7_s1_address),                         //                                hex4_7_s1.address
		.hex4_7_s1_write                                (mm_interconnect_0_hex4_7_s1_write),                           //                                         .write
		.hex4_7_s1_readdata                             (mm_interconnect_0_hex4_7_s1_readdata),                        //                                         .readdata
		.hex4_7_s1_writedata                            (mm_interconnect_0_hex4_7_s1_writedata),                       //                                         .writedata
		.hex4_7_s1_chipselect                           (mm_interconnect_0_hex4_7_s1_chipselect),                      //                                         .chipselect
		.High_Res_Timer_s1_address                      (mm_interconnect_0_high_res_timer_s1_address),                 //                        High_Res_Timer_s1.address
		.High_Res_Timer_s1_write                        (mm_interconnect_0_high_res_timer_s1_write),                   //                                         .write
		.High_Res_Timer_s1_readdata                     (mm_interconnect_0_high_res_timer_s1_readdata),                //                                         .readdata
		.High_Res_Timer_s1_writedata                    (mm_interconnect_0_high_res_timer_s1_writedata),               //                                         .writedata
		.High_Res_Timer_s1_chipselect                   (mm_interconnect_0_high_res_timer_s1_chipselect),              //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.KEYS_s1_address                                (mm_interconnect_0_keys_s1_address),                           //                                  KEYS_s1.address
		.KEYS_s1_write                                  (mm_interconnect_0_keys_s1_write),                             //                                         .write
		.KEYS_s1_readdata                               (mm_interconnect_0_keys_s1_readdata),                          //                                         .readdata
		.KEYS_s1_writedata                              (mm_interconnect_0_keys_s1_writedata),                         //                                         .writedata
		.KEYS_s1_chipselect                             (mm_interconnect_0_keys_s1_chipselect),                        //                                         .chipselect
		.LEDG_s1_address                                (mm_interconnect_0_ledg_s1_address),                           //                                  LEDG_s1.address
		.LEDG_s1_write                                  (mm_interconnect_0_ledg_s1_write),                             //                                         .write
		.LEDG_s1_readdata                               (mm_interconnect_0_ledg_s1_readdata),                          //                                         .readdata
		.LEDG_s1_writedata                              (mm_interconnect_0_ledg_s1_writedata),                         //                                         .writedata
		.LEDG_s1_chipselect                             (mm_interconnect_0_ledg_s1_chipselect),                        //                                         .chipselect
		.ledr_s1_address                                (mm_interconnect_0_ledr_s1_address),                           //                                  ledr_s1.address
		.ledr_s1_write                                  (mm_interconnect_0_ledr_s1_write),                             //                                         .write
		.ledr_s1_readdata                               (mm_interconnect_0_ledr_s1_readdata),                          //                                         .readdata
		.ledr_s1_writedata                              (mm_interconnect_0_ledr_s1_writedata),                         //                                         .writedata
		.ledr_s1_chipselect                             (mm_interconnect_0_ledr_s1_chipselect),                        //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.sbus_decoder_channel_0_s1_address              (mm_interconnect_0_sbus_decoder_channel_0_s1_address),         //                sbus_decoder_channel_0_s1.address
		.sbus_decoder_channel_0_s1_readdata             (mm_interconnect_0_sbus_decoder_channel_0_s1_readdata),        //                                         .readdata
		.sbus_decoder_channel_1_s1_address              (mm_interconnect_0_sbus_decoder_channel_1_s1_address),         //                sbus_decoder_channel_1_s1.address
		.sbus_decoder_channel_1_s1_readdata             (mm_interconnect_0_sbus_decoder_channel_1_s1_readdata),        //                                         .readdata
		.sbus_decoder_channel_10_s1_address             (mm_interconnect_0_sbus_decoder_channel_10_s1_address),        //               sbus_decoder_channel_10_s1.address
		.sbus_decoder_channel_10_s1_readdata            (mm_interconnect_0_sbus_decoder_channel_10_s1_readdata),       //                                         .readdata
		.sbus_decoder_channel_11_s1_address             (mm_interconnect_0_sbus_decoder_channel_11_s1_address),        //               sbus_decoder_channel_11_s1.address
		.sbus_decoder_channel_11_s1_readdata            (mm_interconnect_0_sbus_decoder_channel_11_s1_readdata),       //                                         .readdata
		.sbus_decoder_channel_12_s1_address             (mm_interconnect_0_sbus_decoder_channel_12_s1_address),        //               sbus_decoder_channel_12_s1.address
		.sbus_decoder_channel_12_s1_readdata            (mm_interconnect_0_sbus_decoder_channel_12_s1_readdata),       //                                         .readdata
		.sbus_decoder_channel_13_s1_address             (mm_interconnect_0_sbus_decoder_channel_13_s1_address),        //               sbus_decoder_channel_13_s1.address
		.sbus_decoder_channel_13_s1_readdata            (mm_interconnect_0_sbus_decoder_channel_13_s1_readdata),       //                                         .readdata
		.sbus_decoder_channel_14_s1_address             (mm_interconnect_0_sbus_decoder_channel_14_s1_address),        //               sbus_decoder_channel_14_s1.address
		.sbus_decoder_channel_14_s1_readdata            (mm_interconnect_0_sbus_decoder_channel_14_s1_readdata),       //                                         .readdata
		.sbus_decoder_channel_15_s1_address             (mm_interconnect_0_sbus_decoder_channel_15_s1_address),        //               sbus_decoder_channel_15_s1.address
		.sbus_decoder_channel_15_s1_readdata            (mm_interconnect_0_sbus_decoder_channel_15_s1_readdata),       //                                         .readdata
		.sbus_decoder_channel_2_s1_address              (mm_interconnect_0_sbus_decoder_channel_2_s1_address),         //                sbus_decoder_channel_2_s1.address
		.sbus_decoder_channel_2_s1_readdata             (mm_interconnect_0_sbus_decoder_channel_2_s1_readdata),        //                                         .readdata
		.sbus_decoder_channel_3_s1_address              (mm_interconnect_0_sbus_decoder_channel_3_s1_address),         //                sbus_decoder_channel_3_s1.address
		.sbus_decoder_channel_3_s1_readdata             (mm_interconnect_0_sbus_decoder_channel_3_s1_readdata),        //                                         .readdata
		.sbus_decoder_channel_4_s1_address              (mm_interconnect_0_sbus_decoder_channel_4_s1_address),         //                sbus_decoder_channel_4_s1.address
		.sbus_decoder_channel_4_s1_readdata             (mm_interconnect_0_sbus_decoder_channel_4_s1_readdata),        //                                         .readdata
		.sbus_decoder_channel_5_s1_address              (mm_interconnect_0_sbus_decoder_channel_5_s1_address),         //                sbus_decoder_channel_5_s1.address
		.sbus_decoder_channel_5_s1_readdata             (mm_interconnect_0_sbus_decoder_channel_5_s1_readdata),        //                                         .readdata
		.sbus_decoder_channel_6_s1_address              (mm_interconnect_0_sbus_decoder_channel_6_s1_address),         //                sbus_decoder_channel_6_s1.address
		.sbus_decoder_channel_6_s1_readdata             (mm_interconnect_0_sbus_decoder_channel_6_s1_readdata),        //                                         .readdata
		.sbus_decoder_channel_7_s1_address              (mm_interconnect_0_sbus_decoder_channel_7_s1_address),         //                sbus_decoder_channel_7_s1.address
		.sbus_decoder_channel_7_s1_readdata             (mm_interconnect_0_sbus_decoder_channel_7_s1_readdata),        //                                         .readdata
		.sbus_decoder_channel_8_s1_address              (mm_interconnect_0_sbus_decoder_channel_8_s1_address),         //                sbus_decoder_channel_8_s1.address
		.sbus_decoder_channel_8_s1_readdata             (mm_interconnect_0_sbus_decoder_channel_8_s1_readdata),        //                                         .readdata
		.sbus_decoder_channel_9_s1_address              (mm_interconnect_0_sbus_decoder_channel_9_s1_address),         //                sbus_decoder_channel_9_s1.address
		.sbus_decoder_channel_9_s1_readdata             (mm_interconnect_0_sbus_decoder_channel_9_s1_readdata),        //                                         .readdata
		.sbus_decoder_reg_0_s1_address                  (mm_interconnect_0_sbus_decoder_reg_0_s1_address),             //                    sbus_decoder_reg_0_s1.address
		.sbus_decoder_reg_0_s1_write                    (mm_interconnect_0_sbus_decoder_reg_0_s1_write),               //                                         .write
		.sbus_decoder_reg_0_s1_readdata                 (mm_interconnect_0_sbus_decoder_reg_0_s1_readdata),            //                                         .readdata
		.sbus_decoder_reg_0_s1_writedata                (mm_interconnect_0_sbus_decoder_reg_0_s1_writedata),           //                                         .writedata
		.sbus_decoder_reg_0_s1_chipselect               (mm_interconnect_0_sbus_decoder_reg_0_s1_chipselect),          //                                         .chipselect
		.sbus_decoder_reg_1_s1_address                  (mm_interconnect_0_sbus_decoder_reg_1_s1_address),             //                    sbus_decoder_reg_1_s1.address
		.sbus_decoder_reg_1_s1_write                    (mm_interconnect_0_sbus_decoder_reg_1_s1_write),               //                                         .write
		.sbus_decoder_reg_1_s1_readdata                 (mm_interconnect_0_sbus_decoder_reg_1_s1_readdata),            //                                         .readdata
		.sbus_decoder_reg_1_s1_writedata                (mm_interconnect_0_sbus_decoder_reg_1_s1_writedata),           //                                         .writedata
		.sbus_decoder_reg_1_s1_chipselect               (mm_interconnect_0_sbus_decoder_reg_1_s1_chipselect),          //                                         .chipselect
		.sbus_decoder_reg_10_s1_address                 (mm_interconnect_0_sbus_decoder_reg_10_s1_address),            //                   sbus_decoder_reg_10_s1.address
		.sbus_decoder_reg_10_s1_write                   (mm_interconnect_0_sbus_decoder_reg_10_s1_write),              //                                         .write
		.sbus_decoder_reg_10_s1_readdata                (mm_interconnect_0_sbus_decoder_reg_10_s1_readdata),           //                                         .readdata
		.sbus_decoder_reg_10_s1_writedata               (mm_interconnect_0_sbus_decoder_reg_10_s1_writedata),          //                                         .writedata
		.sbus_decoder_reg_10_s1_chipselect              (mm_interconnect_0_sbus_decoder_reg_10_s1_chipselect),         //                                         .chipselect
		.sbus_decoder_reg_2_s1_address                  (mm_interconnect_0_sbus_decoder_reg_2_s1_address),             //                    sbus_decoder_reg_2_s1.address
		.sbus_decoder_reg_2_s1_write                    (mm_interconnect_0_sbus_decoder_reg_2_s1_write),               //                                         .write
		.sbus_decoder_reg_2_s1_readdata                 (mm_interconnect_0_sbus_decoder_reg_2_s1_readdata),            //                                         .readdata
		.sbus_decoder_reg_2_s1_writedata                (mm_interconnect_0_sbus_decoder_reg_2_s1_writedata),           //                                         .writedata
		.sbus_decoder_reg_2_s1_chipselect               (mm_interconnect_0_sbus_decoder_reg_2_s1_chipselect),          //                                         .chipselect
		.sbus_decoder_reg_3_s1_address                  (mm_interconnect_0_sbus_decoder_reg_3_s1_address),             //                    sbus_decoder_reg_3_s1.address
		.sbus_decoder_reg_3_s1_write                    (mm_interconnect_0_sbus_decoder_reg_3_s1_write),               //                                         .write
		.sbus_decoder_reg_3_s1_readdata                 (mm_interconnect_0_sbus_decoder_reg_3_s1_readdata),            //                                         .readdata
		.sbus_decoder_reg_3_s1_writedata                (mm_interconnect_0_sbus_decoder_reg_3_s1_writedata),           //                                         .writedata
		.sbus_decoder_reg_3_s1_chipselect               (mm_interconnect_0_sbus_decoder_reg_3_s1_chipselect),          //                                         .chipselect
		.sbus_decoder_reg_4_s1_address                  (mm_interconnect_0_sbus_decoder_reg_4_s1_address),             //                    sbus_decoder_reg_4_s1.address
		.sbus_decoder_reg_4_s1_write                    (mm_interconnect_0_sbus_decoder_reg_4_s1_write),               //                                         .write
		.sbus_decoder_reg_4_s1_readdata                 (mm_interconnect_0_sbus_decoder_reg_4_s1_readdata),            //                                         .readdata
		.sbus_decoder_reg_4_s1_writedata                (mm_interconnect_0_sbus_decoder_reg_4_s1_writedata),           //                                         .writedata
		.sbus_decoder_reg_4_s1_chipselect               (mm_interconnect_0_sbus_decoder_reg_4_s1_chipselect),          //                                         .chipselect
		.sbus_decoder_reg_5_s1_address                  (mm_interconnect_0_sbus_decoder_reg_5_s1_address),             //                    sbus_decoder_reg_5_s1.address
		.sbus_decoder_reg_5_s1_write                    (mm_interconnect_0_sbus_decoder_reg_5_s1_write),               //                                         .write
		.sbus_decoder_reg_5_s1_readdata                 (mm_interconnect_0_sbus_decoder_reg_5_s1_readdata),            //                                         .readdata
		.sbus_decoder_reg_5_s1_writedata                (mm_interconnect_0_sbus_decoder_reg_5_s1_writedata),           //                                         .writedata
		.sbus_decoder_reg_5_s1_chipselect               (mm_interconnect_0_sbus_decoder_reg_5_s1_chipselect),          //                                         .chipselect
		.sbus_decoder_reg_6_s1_address                  (mm_interconnect_0_sbus_decoder_reg_6_s1_address),             //                    sbus_decoder_reg_6_s1.address
		.sbus_decoder_reg_6_s1_write                    (mm_interconnect_0_sbus_decoder_reg_6_s1_write),               //                                         .write
		.sbus_decoder_reg_6_s1_readdata                 (mm_interconnect_0_sbus_decoder_reg_6_s1_readdata),            //                                         .readdata
		.sbus_decoder_reg_6_s1_writedata                (mm_interconnect_0_sbus_decoder_reg_6_s1_writedata),           //                                         .writedata
		.sbus_decoder_reg_6_s1_chipselect               (mm_interconnect_0_sbus_decoder_reg_6_s1_chipselect),          //                                         .chipselect
		.sbus_decoder_reg_7_s1_address                  (mm_interconnect_0_sbus_decoder_reg_7_s1_address),             //                    sbus_decoder_reg_7_s1.address
		.sbus_decoder_reg_7_s1_write                    (mm_interconnect_0_sbus_decoder_reg_7_s1_write),               //                                         .write
		.sbus_decoder_reg_7_s1_readdata                 (mm_interconnect_0_sbus_decoder_reg_7_s1_readdata),            //                                         .readdata
		.sbus_decoder_reg_7_s1_writedata                (mm_interconnect_0_sbus_decoder_reg_7_s1_writedata),           //                                         .writedata
		.sbus_decoder_reg_7_s1_chipselect               (mm_interconnect_0_sbus_decoder_reg_7_s1_chipselect),          //                                         .chipselect
		.sbus_decoder_reg_8_s1_address                  (mm_interconnect_0_sbus_decoder_reg_8_s1_address),             //                    sbus_decoder_reg_8_s1.address
		.sbus_decoder_reg_8_s1_write                    (mm_interconnect_0_sbus_decoder_reg_8_s1_write),               //                                         .write
		.sbus_decoder_reg_8_s1_readdata                 (mm_interconnect_0_sbus_decoder_reg_8_s1_readdata),            //                                         .readdata
		.sbus_decoder_reg_8_s1_writedata                (mm_interconnect_0_sbus_decoder_reg_8_s1_writedata),           //                                         .writedata
		.sbus_decoder_reg_8_s1_chipselect               (mm_interconnect_0_sbus_decoder_reg_8_s1_chipselect),          //                                         .chipselect
		.sbus_decoder_reg_9_s1_address                  (mm_interconnect_0_sbus_decoder_reg_9_s1_address),             //                    sbus_decoder_reg_9_s1.address
		.sbus_decoder_reg_9_s1_write                    (mm_interconnect_0_sbus_decoder_reg_9_s1_write),               //                                         .write
		.sbus_decoder_reg_9_s1_readdata                 (mm_interconnect_0_sbus_decoder_reg_9_s1_readdata),            //                                         .readdata
		.sbus_decoder_reg_9_s1_writedata                (mm_interconnect_0_sbus_decoder_reg_9_s1_writedata),           //                                         .writedata
		.sbus_decoder_reg_9_s1_chipselect               (mm_interconnect_0_sbus_decoder_reg_9_s1_chipselect),          //                                         .chipselect
		.sdram_0_s1_address                             (mm_interconnect_0_sdram_0_s1_address),                        //                               sdram_0_s1.address
		.sdram_0_s1_write                               (mm_interconnect_0_sdram_0_s1_write),                          //                                         .write
		.sdram_0_s1_read                                (mm_interconnect_0_sdram_0_s1_read),                           //                                         .read
		.sdram_0_s1_readdata                            (mm_interconnect_0_sdram_0_s1_readdata),                       //                                         .readdata
		.sdram_0_s1_writedata                           (mm_interconnect_0_sdram_0_s1_writedata),                      //                                         .writedata
		.sdram_0_s1_byteenable                          (mm_interconnect_0_sdram_0_s1_byteenable),                     //                                         .byteenable
		.sdram_0_s1_readdatavalid                       (mm_interconnect_0_sdram_0_s1_readdatavalid),                  //                                         .readdatavalid
		.sdram_0_s1_waitrequest                         (mm_interconnect_0_sdram_0_s1_waitrequest),                    //                                         .waitrequest
		.sdram_0_s1_chipselect                          (mm_interconnect_0_sdram_0_s1_chipselect),                     //                                         .chipselect
		.switches0_17_s1_address                        (mm_interconnect_0_switches0_17_s1_address),                   //                          switches0_17_s1.address
		.switches0_17_s1_readdata                       (mm_interconnect_0_switches0_17_s1_readdata),                  //                                         .readdata
		.System_Timer_s1_address                        (mm_interconnect_0_system_timer_s1_address),                   //                          System_Timer_s1.address
		.System_Timer_s1_write                          (mm_interconnect_0_system_timer_s1_write),                     //                                         .write
		.System_Timer_s1_readdata                       (mm_interconnect_0_system_timer_s1_readdata),                  //                                         .readdata
		.System_Timer_s1_writedata                      (mm_interconnect_0_system_timer_s1_writedata),                 //                                         .writedata
		.System_Timer_s1_chipselect                     (mm_interconnect_0_system_timer_s1_chipselect),                //                                         .chipselect
		.uart_0_s1_address                              (mm_interconnect_0_uart_0_s1_address),                         //                                uart_0_s1.address
		.uart_0_s1_write                                (mm_interconnect_0_uart_0_s1_write),                           //                                         .write
		.uart_0_s1_read                                 (mm_interconnect_0_uart_0_s1_read),                            //                                         .read
		.uart_0_s1_readdata                             (mm_interconnect_0_uart_0_s1_readdata),                        //                                         .readdata
		.uart_0_s1_writedata                            (mm_interconnect_0_uart_0_s1_writedata),                       //                                         .writedata
		.uart_0_s1_begintransfer                        (mm_interconnect_0_uart_0_s1_begintransfer),                   //                                         .begintransfer
		.uart_0_s1_chipselect                           (mm_interconnect_0_uart_0_s1_chipselect)                       //                                         .chipselect
	);

	ECE178_nios_20_1_irq_mapper irq_mapper (
		.clk           (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (sys_sdram_pll_0_reset_source_reset), // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (sys_sdram_pll_0_reset_source_reset),     // reset_in1.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
